			----------------------------------------------------------------------------------
			-- Company: 
			-- Engineer: 
			-- 
			-- Create Date:    11:32:59 11/17/2017 
			-- Design Name: 
			-- Module Name:    Memory - Memory 
			-- Project Name: 
			-- Target Devices: 
			-- Tool versions: 
			-- Description: 
			--
			-- Dependencies: 
			--
			-- Revision: 
			-- Revision 0.01 - File Created
			-- Additional Comments: 
			--
			----------------------------------------------------------------------------------
			library IEEE;
			use IEEE.STD_LOGIC_1164.ALL;

			-- Uncomment the following library declaration if using
			-- arithmetic functions with Signed or Unsigned values
			use IEEE.NUMERIC_STD.ALL;

			-- Uncomment the following library declaration if instantiating
			-- any Xilinx primitives in this code.
			--library UNISIM;
			--use UNISIM.VComponents.all;

			entity Memory is
				 Port ( Address : in  STD_LOGIC_VECTOR (28 downto 0);
						  Data_In : in  STD_LOGIC_VECTOR (7 downto 0);
						  Data_Out : out  STD_LOGIC_VECTOR (7 downto 0):= (others => '0');
						  R_W : in  STD_LOGIC_vector (1 downto 0));
			end Memory;

			architecture Memory of Memory is
			type Regs1024x128x8 is array (0 to 2**22-1 ) of std_logic_vector (7 downto 0);
	--		type Regs1024x128x8 is array (2**17-1 downto 0, 2**12-1 downto 0) of std_logic_vector (7 downto 0);
			--signal cache_mem: regs1024x128x8;
			begin
			
				process(Address, Data_In, R_W) --0					1				2				3				4
				variable Memory: regs1024x128x8:=("11010010",	"00100000",	"00000000",	"00010110",	"10000000",		 				--0
				                                  "11001110",	"00000000",	"00000000",	"00000000",	"01000001",		 				--5
				                                  "11001110",	"00000000",	"00000000",	"00000001",	"10000010",		 				--A
				                                  "11001110",	"00000000",	"00000000",	"00010111",	"11000110",	    				--F
															 "00101000",	"00000000",	"00000000",	"00000000",	"00000011",		 				--14
															 "11111110",	"00000000",	"00000000",	"00000000",	"00000000",		 				--19
															 "11111110",	"00000000",	"00000000",	"00000000",	"00000000",		 				--1E
															 "11111110",	"00000000",	"00000000",	"00000000",	"00000000",       			--23
				                                  "00110000",	"00011000",	"00100000",	"00000000",	"00000100",       			--28
				                                  "00011000",	"00000000",	"00100000",	"00000000",	"00000001",       			--2D
				                                  "11111110",	"00000000",	"00000000",	"00000000",	"00000000",       			--32
				                                  "11111110",	"00000000",	"00000000",	"00000000",	"00000000",       			--37
				                                  "00000000",	"00101000",	"10000000",	"00000000",	"00000101",		 				--3C
				                                  "00100000",	"00001000",	"01000000",	"00000000",	"00000000",       			--41
				                                  "10110100",	"01000111",	"11111111",	"11110111",	"01000000",						--46
															 "11111110",	"00000000",	"00000000",	"00000000",	"00000000",						--4B                                                                    --75
															 "11001100",   "00110000", "10100000", "00000000", "00000000",       			--50
															 "11100000",	"00000000",	"00000000",	"00000000",	"00000000",       			--55
															 "00000000",	"00000000",	"00000001",	"01110100", "00000000",       			--5A
															 "00000000",	"00000000",	"00000000",	"00000000", "00000000", others=>X"FF");--5F
				begin                                                                                                
						case R_W is                                                                                     
								when "10" => Data_Out<=Memory(to_integer(unsigned(Address(22 downto 0))));
								when "11" => Memory(to_integer(unsigned(Address(22 downto 0)))):=Data_In;
								when others => null;
						end case;
				end process;
--					when '0' => Data_Out<=Memory(to_integer(unsigned(Address(28 downto 12))),to_integer(unsigned(Address(11 downto 0))));
--					when '1' => Memory(to_integer(unsigned(Address(28 downto 12))),to_integer(unsigned(Address(11 downto 0)))):=Data_In;
			end Memory;
--				variable Memory: regs1024x128x8:=("11010010",	"00100000",	"00000000",	"00010100",	"00000000",		 				--0
--				                                  "11010010",	"00100000",	"00000000",	"00010101",	"01000001",		 				--5
--				                                  "11010010",	"00100000",	"00000000",	"00010110",	"10000010",		 				--A
--				                                  "11010010",	"00100000",	"00000000",	"00010111",	"11000011",	    				--F
--															 "01110010",	"00000000",	"00000000",	"00000000",	"00000100",		 				--14
--															 "11111110",	"00100000",	"00000000",	"00000000",	"00000000",		 				--19
--															 "00101010",	"00000000",	"00000010",	"00100100",	"01000101",		 				--1E
--															 "11111110",	"00100000",	"00000000",	"00000000",	"00000100",       			--23
--				                                  "00110000",	"00000000",	"01000000",	"00000000",	"00000110",       			--28
--				                                  "00000000",	"00010000",	"01100000",	"00000000",	"00000111",       			--2D
--				                                  "00100000",	"00010000",	"01100000",	"00000000",	"00000000",       			--32
--				                                  "11111110",	"00100000",	"00000000",	"00000000",	"00000000",       			--37
--				                                  "11111110",	"00100000",	"00000000",	"00000000",	"00000000",		 				--3C
--				                                  "11111110",	"00100000",	"00000000",	"00000000",	"00000000",       			--41
--				                                  "11111110",	"00100000",	"00000000",	"00000000",	"00000000",       			--46                                                                    --75
--															 "11111110",   "00100000", "00000000", "00000000", "00000000",       			--4B
--															 "00000000",	"00100011",	"11100010",	"11101001",	"00000000",       			--50
--															 "00000000",	"00000000",	"00000110",	"11101100", "00000000",       			--55
--															 "00000000",	"00000000",	"11111000",	"01101000", "00000000",       			--5A
--                                            "00000000",	"00000000",	"00000001",	"01001111", "00000000", others=>X"FF");--5F
